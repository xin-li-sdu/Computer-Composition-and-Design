`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/10/17 19:35:00
// Design Name: 
// Module Name: adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module add_sub(
    input [3:0] a, //��λ�з���������
    input [3:0] b, //��λ�з���������
    input cin, //��λ���Ľ�λ�ź�
    input operator, //�����ӷ����Ǽ����� 0��ʾ�ӷ���1��ʾ����
    output [3:0] result, //������������ʽ 
    output overflow //�����־
); 

    
endmodule
