`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/10/17 19:35:00
// Design Name: 
// Module Name: adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_4(
    input [3:0] a,  // 4λ�޷�����
    input [3:0] b, // 4λ�޷�����
    input cin, // ���λ�����Ľ�λ�ź�
    output [3:0] s, // ��λ�͵Ĳ�����ʽ
    output cf // ��λ��־
);
  
    
endmodule
